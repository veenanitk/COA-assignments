// ROUNAK MODI & VEENA NAGAR//17CO236 & 17C0151//15 october 2018`include "fulladder.v"module fulladder_tb;	reg [0:0] a;	reg [0:0] b;	reg [0:0] c;	wire [0:0] sum;	wire [0:0] carry;fulladder d(.a(a),.b(b),.c(c),.sum(sum),.carry(carry));initial begin	$dumpfile("fulladder.vcd");	$dumpvars(0,fulladder_tb);	$monitor("sum=%b , carry=%b ",sum,carry);	a[0]=0;	b[0]=0;	c[0]=0;	#10  a[0]=0;	     b[0]=1;	     c[0]=1;	#10 $finish;endendmodule	